`timescale 1 ps / 1 ps
module icon_bscan_bufg (
  input  wire        DRCK_LOCAL_I,
  output wire        DRCK_LOCAL_O
  );
  assign DRCK_LOCAL_O = DRCK_LOCAL_I;
endmodule
